module mein

// import r2.pipe
// import zenith391.vgtk3.gtk


pub fn entry(core &R2) {
	hello_world := core.cmd('?e hello world')
	eprintln('hello_world $hello_world')

}
